module DataExt(A,Din,Op,DOut);
input[1:0] A;
input[2:0] Op;
input[31:0] Din;
output[31:0] DOut;
assign DOut=(Op==3'b000)?Din:                        //����չ

            (Op==3'b001&&A==2'b00)?{{24{1'b0}},Din[7:0]}:            //�޷����ֽ�
				(Op==3'b001&&A==2'b01)?{{24{1'b0}},Din[15:8]}:
				(Op==3'b001&&A==2'b10)?{{24{1'b0}},Din[23:16]}:
				(Op==3'b001&&A==2'b11)?{{24{1'b0}},Din[31:24]}:
				
            (Op==3'b010&&A==2'b00)?{{24{Din[7]}},Din[7:0]}:            //�з����ֽ�
				(Op==3'b010&&A==2'b01)?{{24{Din[15]}},Din[15:8]}:
				(Op==3'b010&&A==2'b10)?{{24{Din[23]}},Din[23:16]}:
				(Op==3'b010&&A==2'b11)?{{24{Din[31]}},Din[31:24]}:
				
            (Op==3'b011&&A==2'b00)?{{16{1'b0}},Din[15:0]}:              //�޷��Ű���
				(Op==3'b011&&A==2'b01)?{{16{1'b0}},Din[15:0]}: 
				(Op==3'b011&&A==2'b10)?{{16{1'b0}},Din[31:16]}:	
            (Op==3'b011&&A==2'b11)?{{16{1'b0}},Din[31:16]}:					
				
            (Op==3'b100&&A==2'b10)?{{16{Din[31]}},Din[31:16]}:          //�з��Ű���
				(Op==3'b100&&A==2'b11)?{{16{Din[31]}},Din[31:16]}:   
				(Op==3'b100&&A==2'b01)?{{16{Din[15]}},Din[15:0]}:
				(Op==3'b100&&A==2'b00)?{{16{Din[15]}},Din[15:0]}:0;
				
endmodule
