module comp(ax);


endmodule
