module alu_test;
wire[31:0] result;
wire zero;
ALU ew(1,10,-10,result,zero);
endmodule
